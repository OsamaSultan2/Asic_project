module $_DLATCH_N_ (input D, E, output Q);
    DLL_X1 _TECHMAP_REPLACE_ (.D(D), .GN(E), .Q(Q));
endmodule